library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity PM is
  port(
    addr : in unsigned(9 downto 0);
    data_out : out unsigned(31 downto 0)
  );
end PM;

architecture func of PM is

  constant I_NOP   : unsigned(5 downto 0) := "000000";
  constant I_LD    : unsigned(5 downto 0) := "000001";
  constant I_LDS   : unsigned(5 downto 0) := "000010";
  constant I_LDI   : unsigned(5 downto 0) := "000011";
  constant I_ST    : unsigned(5 downto 0) := "000100";
  constant I_STS   : unsigned(5 downto 0) := "000101";
  constant I_SUBI  : unsigned(5 downto 0) := "000110";
  constant I_LSR   : unsigned(5 downto 0) := "000111";
  constant I_LSL   : unsigned(5 downto 0) := "001000";
  constant I_OR    : unsigned(5 downto 0) := "001001";
  constant I_CMP   : unsigned(5 downto 0) := "001010";
  constant I_CMPI  : unsigned(5 downto 0) := "001011";
  constant I_JMP   : unsigned(5 downto 0) := "001100";
  constant I_BRNE  : unsigned(5 downto 0) := "001101";
  constant I_BREQ  : unsigned(5 downto 0) := "001110";
  constant I_BRMI  : unsigned(5 downto 0) := "001111";
  constant I_BRPL  : unsigned(5 downto 0) := "010000";
  constant I_SUB   : unsigned(5 downto 0) := "010001";
  constant I_ADD   : unsigned(5 downto 0) := "010010";
  constant I_ADDI  : unsigned(5 downto 0) := "010011";
  constant I_INC   : unsigned(5 downto 0) := "010100";
  constant I_DEC   : unsigned(5 downto 0) := "010101";
  constant I_AND   : unsigned(5 downto 0) := "010110";
  constant I_ANDI  : unsigned(5 downto 0) := "010111";
  constant I_ORI   : unsigned(5 downto 0) := "011000";

  constant r0      : unsigned(7 downto 0) := X"00";
  constant r1      : unsigned(7 downto 0) := X"01";
  constant r2      : unsigned(7 downto 0) := X"02";
  constant r3      : unsigned(7 downto 0) := X"03";
  constant r4      : unsigned(7 downto 0) := X"04";
  constant r5      : unsigned(7 downto 0) := X"05";
  constant r6      : unsigned(7 downto 0) := X"06";
  constant r7      : unsigned(7 downto 0) := X"07";
  constant r8      : unsigned(7 downto 0) := X"08";
  constant r9      : unsigned(7 downto 0) := X"09";

  constant audio   : unsigned(9 downto 0) := "0110001100";
  constant key_start : unsigned(9 downto 0) := b"01_1000_1101";
	constant key_2 : unsigned(9 downto 0) := b"01_1000_1110";
	constant DM        : unsigned(9 downto 0) := b"01_1001_0110";

  constant NOP : unsigned(31 downto 0) := X"00000000";

  type PM_t is array(0 to 255) of unsigned(31 downto 0);
  constant PM_c : PM_t := (
--Labels: {'CHORD_HANDLED': 97, 'CHORD_SUCCEEDED': 76, 'OLD_NOTE_SPRITE': 128, 'NEW_NOTE_SPRITE': 150, 'TICK': 122, 'DRAW_TILE_ROW': 2, 'INIT': 0, 'MOVE_BUTTON_INDICATOR': 24, 'DRAW_TILE': 9, 'UPDATE_SCORE': 83, 'NOTE_SPRITE_DECIDED': 156, 'OLD_CHORD': 125, 'NEW_CHORD': 134, 'SET_BUTTON_INDICATOR': 102, 'INDICATOR_DECIDED': 107, 'WAIT0': 43, 'WAIT1': 44, 'WAIT2': 45, 'UPDATE_PREV_INPUT': 96, 'DRAW_TILE_COL': 3, 'EXIT': 169, 'KEEP_AUDIO': 63, 'CHORD_FAILED': 92, 'LOOP': 42}
--Variables: {'c_chord_x': '100', 'c_tile_num_guitar': '2', 'c_tile_num_bg': '1', 'c_chord_dy': '32', 'c_numbers_tile_n': '3', 'c_sprite_num_blank_note': '6', 'a_audio_space': '396', 'a_sprite_n_space_end': '332', 'c_disp_width': '160', 'c_tile_cols': '20', 'a_keyboard_space': '402', 'c_sprite_num_last_note': '5', 'c_strum_y_begin': '96', 'c_guitar_x_end': '13', 'c_strum_y_end': '112', 'a_tile_space_end': '300', 'c_guitar_x_begin': '6', 'c_chord_notes': '5', 'a_keyboard_q': '397', 'a_sprite_x_space_end': '364', 'c_visible_chords': '4', 'a_keyboard_e': '399', 'a_sprite_y_space_begin': '364', 'a_keyboard_w': '398', 'a_keyboard_t': '401', 'c_sprite_num_pressed_note': '7', 'a_keyboard_r': '400', 'a_data_space_begin': '406', 'a_score_tile': '24', 'a_sprite_y_space_end': '396', 'a_tile_space_begin': '0', 'c_tile_rows': '15', 'a_sprite_x_space_begin': '332', 'c_disp_half_height': '60', 'c_note_dx': '12', 'c_disp_height': '120', 'a_sprite_n_space_begin': '300', 'c_strum_y': '104'}
--Registers: {'r_tmp6': 'r20', 'r_score_1': 'r17', 'r_tmp4': 'r27', 'r_tmp5': 'r26', 'r_tmp2': 'r29', 'r_tmp3': 'r28', 'r_tmp0': 'r31', 'r_tmp1': 'r30', 'r_blank_y': 'r2', 'r_blank_x': 'r1', 'r_tile_num': 'r1', 'r_input_space_prev': 'r18', 'r_curr_chord_handled': 'r21', 'r_curr_chord_y': 'r22', 'r_input_space': 'r19', 'r_wait0': 'r10', 'r_wait1': 'r11', 'r_new_note_n': 'r0', 'r_wait2': 'r12', 'r_new_note_y': 'r2', 'r_new_note_x': 'r1', 'r_blank_n': 'r0', 'r_curr_chord_notes': 'r24', 'r_input_qwert': 'r20', 'r_tile_y': 'r3', 'r_curr_chord_addr': 'r25', 'r_tile_x': 'r2', 'r_score_10': 'r16', 'r_tile': 'r0', 'r_curr_chord_audio': 'r23'}
B"000011_00000000_000000000000000000", -- ldi 0b00000000 0 
B"000011_00000011_000000000000000000", -- ldi 0b00000011 0 
B"000011_00000010_000000000000000000", -- ldi 0b00000010 0 
B"000011_00000001_000000000000000001", -- ldi 0b00000001 1 
B"001011_0000000000000010_0000000110", -- cpi 0b00000010 6 
B"001111_00000000000000000000001001", -- brmi 9 
B"001011_0000000000000010_0000001101", -- cpi 0b00000010 13 
B"010000_00000000000000000000001001", -- brpl 9 
B"000011_00000001_000000000000000010", -- ldi 0b00000001 2 
B"000100_00000000_000000010000000000", -- st 0b00000000 0b00000001 
B"010100_00000000_000000000000000000", -- inc 0b00000000 
B"010100_00000010_000000100000000000", -- inc 0b00000010 
B"001011_0000000000000010_0000010100", -- cpi 0b00000010 20 
B"001101_00000000000000000000000011", -- brne 3 
B"010100_00000011_000000110000000000", -- inc 0b00000011 
B"001011_0000000000000011_0000001111", -- cpi 0b00000011 15 
B"001101_00000000000000000000000010", -- brne 2 
B"000011_00000001_000000000001100100", -- ldi 0b00000001 100 
B"000011_00000010_000000000001101000", -- ldi 0b00000010 104 
B"000011_00011111_000000000101001100", -- ldi 0b00011111 332 
B"010011_00011111_00011111_0000000101", -- addi 0b00011111 0b00011111 5 
B"000011_00011110_000000000101101100", -- ldi 0b00011110 364 
B"010011_00011110_00011110_0000000101", -- addi 0b00011110 0b00011110 5 
B"000011_00011101_000000000000000000", -- ldi 0b00011101 0 
B"000100_00011111_000000010000000000", -- st 0b00011111 0b00000001 
B"000100_00011110_000000100000000000", -- st 0b00011110 0b00000010 
B"000110_00000001_00000001_0000001100", -- subi 0b00000001 0b00000001 12 
B"010100_00011111_000111110000000000", -- inc 0b00011111 
B"010100_00011110_000111100000000000", -- inc 0b00011110 
B"010100_00011101_000111010000000000", -- inc 0b00011101 
B"001011_0000000000011101_0000000101", -- cpi 0b00011101 5 
B"001101_00000000000000000000011000", -- brne 24 
B"000011_00011111_000000000000011000", -- ldi 0b00011111 24 
B"000011_00011110_000000000000000011", -- ldi 0b00011110 3 
B"000100_00011111_000111100000000000", -- st 0b00011111 0b00011110 
B"010101_00011111_000111110000000000", -- dec 0b00011111 
B"000100_00011111_000111100000000000", -- st 0b00011111 0b00011110 
B"000011_00010110_000000000001111000", -- ldi 0b00010110 120 
B"000011_00011001_000000000110010110", -- ldi 0b00011001 406 
B"000011_00010101_000000000000000000", -- ldi 0b00010101 0 
B"000011_00010001_000000000000000000", -- ldi 0b00010001 0 
B"000011_00010000_000000000000000000", -- ldi 0b00010000 0 
B"000011_00001010_000000000000001111", -- ldi 0b00001010 15 
B"000011_00001011_000000000111111111", -- ldi 0b00001011 511 
B"000011_00001100_000000000000000001", -- ldi 0b00001100 1 
B"000010_00010100_000000000110001101", -- lds 0b00010100 397 
B"001000_00010100_00010100_0000000001", -- lsl 0b00010100 1 
B"000010_00011111_000000000110001110", -- lds 0b00011111 398 
B"001001_00010100_00010100_0001111100", -- or 0b00010100 0b00010100 0b00011111 
B"001000_00010100_00010100_0000000001", -- lsl 0b00010100 1 
B"000010_00011111_000000000110001111", -- lds 0b00011111 399 
B"001001_00010100_00010100_0001111100", -- or 0b00010100 0b00010100 0b00011111 
B"001000_00010100_00010100_0000000001", -- lsl 0b00010100 1 
B"000010_00011111_000000000110010000", -- lds 0b00011111 400 
B"001001_00010100_00010100_0001111100", -- or 0b00010100 0b00010100 0b00011111 
B"001000_00010100_00010100_0000000001", -- lsl 0b00010100 1 
B"000010_00011111_000000000110010001", -- lds 0b00011111 401 
B"001001_00010100_00010100_0001111100", -- or 0b00010100 0b00010100 0b00011111 
B"000010_00010011_000000000110010010", -- lds 0b00010011 402 
B"001011_0000000000010110_0000111100", -- cpi 0b00010110 60 
B"001101_00000000000000000000111111", -- brne 63 
B"000011_00011111_000000000000000000", -- ldi 0b00011111 0 
B"000101_0000000000011111_0110001100", -- sts 396 0b00011111 
B"001011_0000000000010101_0000000000", -- cpi 0b00010101 0 
B"001101_00000000000000000001100001", -- brne 97 
B"001011_0000000000010011_0000000001", -- cpi 0b00010011 1 
B"001101_00000000000000000001100000", -- brne 96 
B"001011_0000000000010010_0000000000", -- cpi 0b00010010 0 
B"001101_00000000000000000001100001", -- brne 97 
B"000011_00010010_000000000000000001", -- ldi 0b00010010 1 
B"001011_0000000000010110_0001100000", -- cpi 0b00010110 96 
B"001111_00000000000000000001011100", -- brmi 92 
B"001011_0000000000010110_0001110000", -- cpi 0b00010110 112 
B"010000_00000000000000000001011100", -- brpl 92 
B"001010_0000000000011000_0001010000", -- cp 0b00011000 0b00010100 
B"001101_00000000000000000001011100", -- brne 92 
B"000011_00010101_000000000000000001", -- ldi 0b00010101 1 
B"000101_0000000000010111_0110001100", -- sts 396 0b00010111 
B"010100_00010001_000100010000000000", -- inc 0b00010001 
B"001011_0000000000010001_0000001010", -- cpi 0b00010001 10 
B"001101_00000000000000000001010011", -- brne 83 
B"000011_00010001_000000000000000000", -- ldi 0b00010001 0 
B"010100_00010000_000100000000000000", -- inc 0b00010000 
B"000011_00011111_000000000000011000", -- ldi 0b00011111 24 
B"000011_00011110_000000000000000011", -- ldi 0b00011110 3 
B"010010_00011110_00011110_0001000100", -- add 0b00011110 0b00011110 0b00010001 
B"000100_00011111_000111100000000000", -- st 0b00011111 0b00011110 
B"010101_00011111_000111110000000000", -- dec 0b00011111 
B"000011_00011110_000000000000000011", -- ldi 0b00011110 3 
B"010010_00011110_00011110_0001000000", -- add 0b00011110 0b00011110 0b00010000 
B"000100_00011111_000111100000000000", -- st 0b00011111 0b00011110 
B"001100_00000000000000000001100001", -- jmp 97 
B"000011_00010101_000000000000000001", -- ldi 0b00010101 1 
B"000011_00011111_000000000000000000", -- ldi 0b00011111 0 
B"000101_0000000000011111_0110001100", -- sts 396 0b00011111 
B"001100_00000000000000000001100001", -- jmp 97 
B"000011_00010010_000000000000000000", -- ldi 0b00010010 0 
B"000011_00011111_000000000100101100", -- ldi 0b00011111 300 
B"010011_00011111_00011111_0000000101", -- addi 0b00011111 0b00011111 5 
B"000011_00011110_000000000000000000", -- ldi 0b00011110 0 
B"000011_00011101_000000000000000000", -- ldi 0b00011101 0 
B"001001_00011101_00011101_0001010000", -- or 0b00011101 0b00011101 0b00010100 
B"000011_00000000_000000000000000110", -- ldi 0b00000000 6 
B"010111_00011100_00011101_0000000001", -- andi 0b00011100 0b00011101 1 
B"001011_0000000000011100_0000000001", -- cpi 0b00011100 1 
B"001101_00000000000000000001101011", -- brne 107 
B"000011_00000000_000000000000000111", -- ldi 0b00000000 7 
B"000100_00011111_000000000000000000", -- st 0b00011111 0b00000000 
B"010100_00011111_000111110000000000", -- inc 0b00011111 
B"000111_00011101_00011101_0000000001", -- lsr 0b00011101 1 
B"010100_00011110_000111100000000000", -- inc 0b00011110 
B"001011_0000000000011110_0000000101", -- cpi 0b00011110 5 
B"001101_00000000000000000001100110", -- brne 102 
B"010101_00001100_000011000000000000", -- dec 0b00001100 
B"001011_0000000000001100_0000000000", -- cpi 0b00001100 0 
B"001101_00000000000000000000101101", -- brne 45 
B"010101_00001011_000010110000000000", -- dec 0b00001011 
B"001011_0000000000001011_0000000000", -- cpi 0b00001011 0 
B"001101_00000000000000000000101100", -- brne 44 
B"010101_00001010_000010100000000000", -- dec 0b00001010 
B"001011_0000000000001010_0000000000", -- cpi 0b00001010 0 
B"001101_00000000000000000000101011", -- brne 43 
B"001011_0000000000010110_0001111000", -- cpi 0b00010110 120 
B"001110_00000000000000000010000110", -- breq 134 
B"001100_00000000000000000001111101", -- jmp 125 
B"010100_00010110_000101100000000000", -- inc 0b00010110 
B"000011_00011111_000000000101101100", -- ldi 0b00011111 364 
B"000011_00011110_000000000000000000", -- ldi 0b00011110 0 
B"000100_00011111_000101100000000000", -- st 0b00011111 0b00010110 
B"010100_00011111_000111110000000000", -- inc 0b00011111 
B"010100_00011110_000111100000000000", -- inc 0b00011110 
B"001011_0000000000011110_0000000101", -- cpi 0b00011110 5 
B"001101_00000000000000000010000000", -- brne 128 
B"001100_00000000000000000000101010", -- jmp 42 
B"000001_00011000_000110010000000000", -- ld 0b00011000 0b00011001 
B"001011_0000000000011000_1111111111", -- cpi 0b00011000 1023 
B"001110_00000000000000000010101001", -- breq 169 
B"000111_00011000_00011000_0000000011", -- lsr 0b00011000 3 
B"000001_00010111_000110010000000000", -- ld 0b00010111 0b00011001 
B"000011_00010110_000000000000000000", -- ldi 0b00010110 0 
B"000011_00010101_000000000000000000", -- ldi 0b00010101 0 
B"000011_00000000_000000000000000101", -- ldi 0b00000000 5 
B"000011_00000001_000000000001100100", -- ldi 0b00000001 100 
B"000011_00000010_000000000000000000", -- ldi 0b00000010 0 
B"000011_00011111_000000000100101100", -- ldi 0b00011111 300 
B"000011_00011110_000000000101001100", -- ldi 0b00011110 332 
B"000011_00011101_000000000101101100", -- ldi 0b00011101 364 
B"000011_00011100_000000000000000000", -- ldi 0b00011100 0 
B"000011_00011010_000000000000000000", -- ldi 0b00011010 0 
B"001001_00011010_00011000_0001101000", -- or 0b00011010 0b00011000 0b00011010 
B"000011_00010100_000000000000000000", -- ldi 0b00010100 0 
B"000100_00011111_000101000000000000", -- st 0b00011111 0b00010100 
B"010111_00011011_00011010_0000000001", -- andi 0b00011011 0b00011010 1 
B"001011_0000000000011011_0000000001", -- cpi 0b00011011 1 
B"001101_00000000000000000010011100", -- brne 156 
B"000100_00011111_000000000000000000", -- st 0b00011111 0b00000000 
B"000100_00011110_000000010000000000", -- st 0b00011110 0b00000001 
B"000100_00011101_000000100000000000", -- st 0b00011101 0b00000010 
B"000110_00000001_00000001_0000001100", -- subi 0b00000001 0b00000001 12 
B"010101_00000000_000000000000000000", -- dec 0b00000000 
B"010100_00011111_000111110000000000", -- inc 0b00011111 
B"010100_00011110_000111100000000000", -- inc 0b00011110 
B"010100_00011101_000111010000000000", -- inc 0b00011101 
B"000111_00011010_00011010_0000000001", -- lsr 0b00011010 1 
B"010100_00011100_000111000000000000", -- inc 0b00011100 
B"001011_0000000000011100_0000000101", -- cpi 0b00011100 5 
B"001101_00000000000000000010010110", -- brne 150 
B"010100_00011001_000110010000000000", -- inc 0b00011001 
B"001100_00000000000000000000101010", -- jmp 42 
B"001100_00000000000000000010101001", -- jmp 169 
    others => (others => '0')
    );

begin
  data_out <= PM_c(to_integer(addr));

end architecture;
