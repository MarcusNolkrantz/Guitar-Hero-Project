x"00",x"00",x"e0",x"e0",x"e0",x"e0",x"00",x"00",
x"00",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"00",
x"e0",x"e0",x"e0",x"ff",x"ff",x"e0",x"e0",x"e0",
x"e0",x"e0",x"e0",x"ff",x"ff",x"e0",x"e0",x"e0",
x"e0",x"e0",x"e0",x"9f",x"9f",x"e0",x"e0",x"e0",
x"80",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"80",
x"00",x"80",x"e0",x"e0",x"e0",x"e0",x"80",x"00",
x"00",x"00",x"80",x"80",x"80",x"80",x"00",x"00",
x"00",x"00",x"78",x"78",x"78",x"78",x"00",x"00",
x"00",x"78",x"78",x"78",x"78",x"78",x"78",x"00",
x"78",x"78",x"78",x"ff",x"ff",x"78",x"78",x"78",
x"78",x"78",x"78",x"ff",x"ff",x"78",x"78",x"78",
x"78",x"78",x"78",x"9f",x"9f",x"78",x"78",x"78",
x"10",x"78",x"78",x"78",x"78",x"78",x"78",x"10",
x"00",x"10",x"78",x"78",x"78",x"78",x"10",x"00",
x"00",x"00",x"10",x"10",x"10",x"10",x"00",x"00",
x"00",x"00",x"fc",x"fc",x"fc",x"fc",x"00",x"00",
x"00",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"00",
x"fc",x"fc",x"fc",x"ff",x"ff",x"fc",x"fc",x"fc",
x"fc",x"fc",x"fc",x"ff",x"ff",x"fc",x"fc",x"fc",
x"fc",x"fc",x"fc",x"9f",x"9f",x"fc",x"fc",x"fc",
x"f4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f4",
x"00",x"f4",x"fc",x"fc",x"fc",x"fc",x"f4",x"00",
x"00",x"00",x"f4",x"f4",x"f4",x"f4",x"00",x"00",
x"00",x"00",x"07",x"07",x"07",x"07",x"00",x"00",
x"00",x"07",x"07",x"07",x"07",x"07",x"07",x"00",
x"07",x"07",x"07",x"ff",x"ff",x"07",x"07",x"07",
x"07",x"07",x"07",x"ff",x"ff",x"07",x"07",x"07",
x"07",x"07",x"07",x"9f",x"9f",x"07",x"07",x"07",
x"01",x"07",x"07",x"07",x"07",x"07",x"07",x"01",
x"00",x"01",x"07",x"07",x"07",x"07",x"01",x"00",
x"00",x"00",x"01",x"01",x"01",x"01",x"00",x"00",
x"00",x"00",x"f0",x"f0",x"f0",x"f0",x"00",x"00",
x"00",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"00",
x"f0",x"f0",x"f0",x"ff",x"ff",x"f0",x"f0",x"f0",
x"f0",x"f0",x"f0",x"ff",x"ff",x"f0",x"f0",x"f0",
x"f0",x"f0",x"f0",x"9f",x"9f",x"f0",x"f0",x"f0",
x"b0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"b0",
x"00",x"b0",x"f0",x"f0",x"f0",x"f0",x"b0",x"00",
x"00",x"00",x"b0",x"b0",x"b0",x"b0",x"00",x"00",
