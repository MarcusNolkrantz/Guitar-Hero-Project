x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"0f",x"00",x"00",x"00",x"00",
x"00",x"00",x"0f",x"0f",x"0f",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"0f",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"0f",x"0f",x"00",x"00",
x"00",x"00",x"00",x"0f",x"00",x"0f",x"00",x"00",
x"00",x"00",x"0f",x"0f",x"0f",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"0f",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
