x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",
x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",
x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",
x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",
x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",
x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",
x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",
x"97",x"97",x"97",x"97",x"97",x"97",x"97",x"97",
