x"00",x"04",x"04",x"04",x"04",x"04",x"04",x"00",
x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",
x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",
x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",
x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",
x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",
x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",
x"00",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"00",
