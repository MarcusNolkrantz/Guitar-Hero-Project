x"00",x"00",x"97",x"97",x"97",x"97",x"00",x"00",
x"00",x"97",x"04",x"04",x"04",x"04",x"97",x"00",
x"97",x"04",x"00",x"00",x"00",x"00",x"04",x"97",
x"97",x"00",x"00",x"00",x"00",x"00",x"00",x"97",
x"97",x"00",x"00",x"00",x"00",x"00",x"00",x"97",
x"04",x"97",x"00",x"00",x"00",x"00",x"97",x"04",
x"00",x"04",x"97",x"97",x"97",x"97",x"04",x"00",
x"00",x"00",x"04",x"04",x"04",x"04",x"00",x"00",
