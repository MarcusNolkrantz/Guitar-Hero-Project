x"0f",x"02",x"0a",x"0a",x"0f",x"0a",x"0a",x"02",
x"02",x"0a",x"02",x"0a",x"02",x"0a",x"02",x"0f",
x"0a",x"00",x"00",x"02",x"0a",x"00",x"00",x"0f",
x"0a",x"00",x"00",x"0a",x"02",x"00",x"00",x"0a",
x"02",x"0a",x"0a",x"00",x"00",x"0f",x"02",x"02",
x"0a",x"02",x"00",x"00",x"00",x"00",x"0a",x"0f",
x"0f",x"02",x"00",x"00",x"00",x"00",x"0a",x"02",
x"0a",x"0a",x"00",x"0a",x"0f",x"00",x"02",x"0a",
x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",
x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",
x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",
x"00",x"0f",x"db",x"db",x"db",x"db",x"0f",x"00",
x"db",x"db",x"cf",x"cf",x"cf",x"cf",x"db",x"db",
x"db",x"db",x"c7",x"cf",x"cf",x"c7",x"db",x"db",
x"db",x"db",x"cf",x"cf",x"cf",x"cf",x"db",x"db",
x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
