library ieee;
use ieee.std_logic_1164.ALL;            -- basic IEEE library
use ieee.numeric_std.ALL;               -- IEEE library for the unsigned type

entity DM is
  port (
    clk         : in  std_logic;
    rst         : in  std_logic;
    we          : in  std_logic;
    addr_read   : in  unsigned(9 downto 0);
    data_read   : out std_logic_vector(15 downto 0);
    addr_write  : in  unsigned(9 downto 0);
    data_write  : in  std_logic_vector(15 downto 0)
  );
end entity;

architecture behaviour of DM is

  type DM_t is array (0 to 127) of std_logic_vector(15 downto 0);
  signal DM_content : DM_t := (
    -- blinka lilla stjärna
    "0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000100111",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000001000110",
"0000000010000100",
"0000000000000000",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000100111",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000001000110",
"0000000010000100",
"0000000000000000",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000100111",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000001000110",
"0000000010000100",
"0000000000000000",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000100111",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000001000110",
"0000000010000100",
"0000000000000000",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000100111",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000001000110",
"0000000010000100",
"0000000000000000",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000100111",
"0000000010000100",
"0000000001000110",
"0000000000100111",
"0000000000000000",
"0000000001000110",
"0000000010000100",
"0000000000000000",
"0000000000000000",
    others => (others => '0'))
;

begin
  process(clk) begin
    if rising_edge(clk) then
      if we = '1' then    
          DM_content(to_integer(addr_write)) <= data_write;
	end if;	
	data_read <= DM_content(to_integer(addr_read));
    end if;
  end process;
end architecture;
